** sch_path: /home/edney_freitas/Tutorial/inverter_tutorial/xschem/inverter.sch
.subckt inverter VDD Vout Vin VSS
*.ipin Vin
*.iopin VDD
*.iopin Vout
*.iopin VSS
XM1 Vout Vin VSS VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM2 Vout Vin VDD VDD sg13_lv_pmos w=3u l=0.13u ng=1 m=1
.ends
.end
