* Extracted by KLayout with SG13G2 LVS runset on : 29/01/2026 08:25

.SUBCKT inverter
M$1 \$1 \$3 \$2 \$1 sg13_lv_nmos L=0.13u W=1u AS=0.34p AD=0.34p PS=2.68u
+ PD=2.68u
M$2 \$4 \$3 \$2 \$4 sg13_lv_pmos L=0.13u W=3u AS=1.02p AD=1.02p PS=6.68u
+ PD=6.68u
.ENDS inverter
