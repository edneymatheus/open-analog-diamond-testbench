** sch_path: /home/jsmoya07/Documents/inverter_tutorial/xschem/inverter_tb.sch
**.subckt inverter_tb
x1 VDD Vout Vin VSS inverter
C1 Vout VSS 100f m=1
V1 VSS GND 0
V2 VDD VSS 1.5
V3 Vin VSS 1.5
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt



.dc V3 0 1.5 0.01
.save all


**** end user architecture code
**.ends

* expanding   symbol:  /home/jsmoya07/Documents/inverter_tutorial/xschem/inverter.sym # of pins=4
** sym_path: /home/jsmoya07/Documents/inverter_tutorial/xschem/inverter.sym
** sch_path: /home/jsmoya07/Documents/inverter_tutorial/xschem/inverter.sch
.subckt inverter VDD Vout Vin VSS
*.ipin Vin
*.iopin VDD
*.iopin Vout
*.iopin VSS
XM1 Vout Vin VSS VSS sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM2 Vout Vin VDD VDD sg13_lv_pmos w=3u l=0.13u ng=1 m=1
.ends

.GLOBAL GND
.end
